/**
 *  Non-linear function Fc enumerator
 *  NLF takes 5 inputs and produces a single output.
 *  fn=0xEC57E80A
 *  This enumerator reverses that and takes a single
 *  input bit to enumerator all states that produce
 *  that bit.
 * 
 *  Elliot Buller
 *  2022
 */

module FcEnum
  (
   input              CLK,
   input              RESETn,
   input              BIT,
   output logic [4:0] OUTPUT
   );
   

endmodule // FcEnum
